// sdram.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module sdram (
		input  wire        clk_clk,                 //       clk.clk
		input  wire        reset_reset,             //     reset.reset
		output wire        sdr_clk_clk,             //   sdr_clk.clk
		input  wire [24:0] sdr_slave_address,       // sdr_slave.address
		input  wire [1:0]  sdr_slave_byteenable_n,  //          .byteenable_n
		input  wire        sdr_slave_chipselect,    //          .chipselect
		input  wire [15:0] sdr_slave_writedata,     //          .writedata
		input  wire        sdr_slave_read_n,        //          .read_n
		input  wire        sdr_slave_write_n,       //          .write_n
		output wire [15:0] sdr_slave_readdata,      //          .readdata
		output wire        sdr_slave_readdatavalid, //          .readdatavalid
		output wire        sdr_slave_waitrequest,   //          .waitrequest
		output wire [12:0] sdr_wire_addr,           //  sdr_wire.addr
		output wire [1:0]  sdr_wire_ba,             //          .ba
		output wire        sdr_wire_cas_n,          //          .cas_n
		output wire        sdr_wire_cke,            //          .cke
		output wire        sdr_wire_cs_n,           //          .cs_n
		inout  wire [15:0] sdr_wire_dq,             //          .dq
		output wire [1:0]  sdr_wire_dqm,            //          .dqm
		output wire        sdr_wire_ras_n,          //          .ras_n
		output wire        sdr_wire_we_n            //          .we_n
	);

	wire    sys_sdram_pll_sys_clk_clk;        // sys_sdram_pll:sys_clk_clk -> [rst_controller:clk, sdram_control:clk]
	wire    rst_controller_reset_out_reset;   // rst_controller:reset_out -> sdram_control:reset_n
	wire    sys_sdram_pll_reset_source_reset; // sys_sdram_pll:reset_source_reset -> rst_controller:reset_in0

	sdram_sdram_control sdram_control (
		.clk            (sys_sdram_pll_sys_clk_clk),       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset), // reset.reset_n
		.az_addr        (sdr_slave_address),               //    s1.address
		.az_be_n        (sdr_slave_byteenable_n),          //      .byteenable_n
		.az_cs          (sdr_slave_chipselect),            //      .chipselect
		.az_data        (sdr_slave_writedata),             //      .writedata
		.az_rd_n        (sdr_slave_read_n),                //      .read_n
		.az_wr_n        (sdr_slave_write_n),               //      .write_n
		.za_data        (sdr_slave_readdata),              //      .readdata
		.za_valid       (sdr_slave_readdatavalid),         //      .readdatavalid
		.za_waitrequest (sdr_slave_waitrequest),           //      .waitrequest
		.zs_addr        (sdr_wire_addr),                   //  wire.export
		.zs_ba          (sdr_wire_ba),                     //      .export
		.zs_cas_n       (sdr_wire_cas_n),                  //      .export
		.zs_cke         (sdr_wire_cke),                    //      .export
		.zs_cs_n        (sdr_wire_cs_n),                   //      .export
		.zs_dq          (sdr_wire_dq),                     //      .export
		.zs_dqm         (sdr_wire_dqm),                    //      .export
		.zs_ras_n       (sdr_wire_ras_n),                  //      .export
		.zs_we_n        (sdr_wire_we_n)                    //      .export
	);

	sdram_sys_sdram_pll sys_sdram_pll (
		.ref_clk_clk        (clk_clk),                          //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                      //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdr_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_reset_source_reset)  // reset_source.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_sdram_pll_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_in1      (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

endmodule
